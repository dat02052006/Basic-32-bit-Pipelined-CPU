library verilog;
use verilog.vl_types.all;
entity CLA32_vlg_check_tst is
    port(
        Sum             : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end CLA32_vlg_check_tst;
