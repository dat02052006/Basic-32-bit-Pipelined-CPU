library verilog;
use verilog.vl_types.all;
entity CLA32_vlg_vec_tst is
end CLA32_vlg_vec_tst;
