library verilog;
use verilog.vl_types.all;
entity bit_slice_vlg_vec_tst is
end bit_slice_vlg_vec_tst;
