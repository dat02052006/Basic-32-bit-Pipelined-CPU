library verilog;
use verilog.vl_types.all;
entity FowardingUnit_vlg_sample_tst is
    port(
        EX_MEM_Rd       : in     vl_logic_vector(4 downto 0);
        EX_MEM_RegWrite : in     vl_logic;
        ID_EX_Rs        : in     vl_logic_vector(4 downto 0);
        ID_EX_Rt        : in     vl_logic_vector(4 downto 0);
        MEM_WB_Rd       : in     vl_logic_vector(4 downto 0);
        MEM_WB_RegWrite : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end FowardingUnit_vlg_sample_tst;
