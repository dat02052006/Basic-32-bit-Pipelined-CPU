library verilog;
use verilog.vl_types.all;
entity CPU_pipeline_vlg_vec_tst is
end CPU_pipeline_vlg_vec_tst;
