library verilog;
use verilog.vl_types.all;
entity FowardingUnit_vlg_vec_tst is
end FowardingUnit_vlg_vec_tst;
