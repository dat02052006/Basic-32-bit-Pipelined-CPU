library verilog;
use verilog.vl_types.all;
entity AL_vlg_vec_tst is
end AL_vlg_vec_tst;
