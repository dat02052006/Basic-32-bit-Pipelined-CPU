library verilog;
use verilog.vl_types.all;
entity Registers_vlg_vec_tst is
end Registers_vlg_vec_tst;
