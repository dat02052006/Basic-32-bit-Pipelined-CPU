library verilog;
use verilog.vl_types.all;
entity RFC32x32_vlg_vec_tst is
end RFC32x32_vlg_vec_tst;
