library verilog;
use verilog.vl_types.all;
entity add4pg_vlg_vec_tst is
end add4pg_vlg_vec_tst;
