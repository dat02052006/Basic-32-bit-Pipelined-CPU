library verilog;
use verilog.vl_types.all;
entity Add4_vlg_vec_tst is
end Add4_vlg_vec_tst;
